module uart_top #(parameter clk_freq = 1000000, parameter baud_rate = 9600)(
    input clk,rst, 
    input rx,
    input [7:0] dintx,
    input newd,
    output tx, 
    output [7:0] doutrx,
    output donetx,
    output donerx
    );
    
    uarttx #(clk_freq, baud_rate) utx (clk, rst, newd, dintx, tx, donetx);   
 
    uartrx #(clk_freq, baud_rate) rtx (clk, rst, rx, donerx, doutrx);    
    
endmodule
